module verification_wrapper(
 input  a0x0_0, a1x0_0, a2x0_0, a3x0_0, a0x1_0, a1x1_0, a2x1_0, a3x1_0, a0x2_0, a1x2_0, a2x2_0, a3x2_0, a0x3_0, a1x3_0, a2x3_0, a3x3_0, a0x4_0, a1x4_0, a2x4_0, a3x4_0, a0x5_0, a1x5_0, a2x5_0, a3x5_0, a0x6_0, a1x6_0, a2x6_0, a3x6_0, a0x7_0, a1x7_0, a2x7_0, a3x7_0,
 input  a0x0_1, a1x0_1, a2x0_1, a3x0_1, a0x1_1, a1x1_1, a2x1_1, a3x1_1, a0x2_1, a1x2_1, a2x2_1, a3x2_1, a0x3_1, a1x3_1, a2x3_1, a3x3_1, a0x4_1, a1x4_1, a2x4_1, a3x4_1, a0x5_1, a1x5_1, a2x5_1, a3x5_1, a0x6_1, a1x6_1, a2x6_1, a3x6_1, a0x7_1, a1x7_1, a2x7_1, a3x7_1,
 input  m0, m1, 
 output b0x0, b1x0, b2x0, b3x0, b0x1, b1x1, b2x1, b3x1, b0x2, b1x2, b2x2, b3x2, b0x3, b1x3, b2x3, b3x3, b0x4, b1x4, b2x4, b3x4, b0x5, b1x5, b2x5, b3x5, b0x6, b1x6, b2x6, b3x6, b0x7, b1x7, b2x7, b3x7);

      // Ensure mask encoding and relation as we assume
      //a0      
      assign a0r0 = (a0x0_0 ^ m1) ^ a0x0_1;      // 2
      assign a0r1 = (a0x1_0 ^ m0 ^ m1) ^ a0x1_1; // 3 
      assign a0r2 = (a0x2_0 ^ m0 ^ m1) ^ a0x2_1; // 3 
      assign a0r3 = (a0x3_0 ^ m0) ^ a0x3_1;      // 1 
      assign a0r4 = (a0x4_0 ^ m0) ^ a0x4_1;      // 1 
      assign a0r5 = (a0x5_0 ^ m1) ^ a0x5_1;      // 2 
      assign a0r6 = (a0x6_0 ^ m0) ^ a0x6_1;      // 1 
      assign a0r7 = (a0x7_0 ^ m1) ^ a0x7_1;      // 2   
      //a1      
      assign a1r0 = (a1x0_0 ^ m1) ^ a1x0_1;      // 2
      assign a1r1 = (a1x1_0 ^ m0 ^ m1) ^ a1x1_1; // 3 
      assign a1r2 = (a1x2_0 ^ m0 ^ m1) ^ a1x2_1; // 3 
      assign a1r3 = (a1x3_0 ^ m0) ^ a1x3_1;      // 1 
      assign a1r4 = (a1x4_0 ^ m0) ^ a1x4_1;      // 1 
      assign a1r5 = (a1x5_0 ^ m1) ^ a1x5_1;      // 2 
      assign a1r6 = (a1x6_0 ^ m0) ^ a1x6_1;      // 1 
      assign a1r7 = (a1x7_0 ^ m1) ^ a1x7_1;      // 2   
      //a2      
      assign a2r0 = (a2x0_0 ^ m1) ^ a2x0_1;      // 2
      assign a2r1 = (a2x1_0 ^ m0 ^ m1) ^ a2x1_1; // 3 
      assign a2r2 = (a2x2_0 ^ m0 ^ m1) ^ a2x2_1; // 3 
      assign a2r3 = (a2x3_0 ^ m0) ^ a2x3_1;      // 1 
      assign a2r4 = (a2x4_0 ^ m0) ^ a2x4_1;      // 1 
      assign a2r5 = (a2x5_0 ^ m1) ^ a2x5_1;      // 2 
      assign a2r6 = (a2x6_0 ^ m0) ^ a2x6_1;      // 1 
      assign a2r7 = (a2x7_0 ^ m1) ^ a2x7_1;      // 2   
      //a3      
      assign a3r0 = (a3x0_0 ^ m1) ^ a3x0_1;      // 2
      assign a3r1 = (a3x1_0 ^ m0 ^ m1) ^ a3x1_1; // 3 
      assign a3r2 = (a3x2_0 ^ m0 ^ m1) ^ a3x2_1; // 3 
      assign a3r3 = (a3x3_0 ^ m0) ^ a3x3_1;      // 1 
      assign a3r4 = (a3x4_0 ^ m0) ^ a3x4_1;      // 1 
      assign a3r5 = (a3x5_0 ^ m1) ^ a3x5_1;      // 2 
      assign a3r6 = (a3x6_0 ^ m0) ^ a3x6_1;      // 1 
      assign a3r7 = (a3x7_0 ^ m1) ^ a3x7_1;      // 2   
      
      // DUV
     mixcolumns mixcolumns_ins(a0r0, a1r0, a2r0, a3r0, a0r1, a1r1, a2r1, a3r1, a0r2, a1r2, a2r2, a3r2, a0r3, a1r3, a2r3, a3r3, a0r4, a1r4, a2r4, a3r4, a0r5, a1r5, a2r5, a3r5, a0r6, a1r6, a2r6, a3r6, a0r7, a1r7, a2r7, a3r7, m0, m1, 
		               b0x0, b1x0, b2x0, b3x0, b0x1, b1x1, b2x1, b3x1, b0x2, b1x2, b2x2, b3x2, b0x3, b1x3, b2x3, b3x3, b0x4, b1x4, b2x4, b3x4, b0x5, b1x5, b2x5, b3x5, b0x6, b1x6, b2x6, b3x6, b0x7, b1x7, b2x7, b3x7);

        
endmodule

/* MixColumns (automatically created) */
module mixcolumns(
	              input  a0x0, a1x0, a2x0, a3x0, a0x1, a1x1, a2x1, a3x1, a0x2, a1x2, a2x2, a3x2, a0x3, a1x3, a2x3, a3x3, a0x4, a1x4, a2x4, a3x4, a0x5, a1x5, a2x5, a3x5, a0x6, a1x6, a2x6, a3x6, a0x7, a1x7, a2x7, a3x7, MASK1, MASK2, 
		          output b0x0, b1x0, b2x0, b3x0, b0x1, b1x1, b2x1, b3x1, b0x2, b1x2, b2x2, b3x2, b0x3, b1x3, b2x3, b3x3, b0x4, b1x4, b2x4, b3x4, b0x5, b1x5, b2x5, b3x5, b0x6, b1x6, b2x6, b3x6, b0x7, b1x7, b2x7, b3x7);
   assign ha0x0_0 = a0x0 ^ MASK1; 
   assign ha0x0_1 = MASK1 ^ MASK2;
   assign a0_mul_2x0_0 = a0x7; 
   assign a0_mul_2x0_1 = MASK2;
   assign a0_mul_2x1_0 = ha0x0_0 ^ a0x7; 
   assign a0_mul_2x1_1 = MASK1;
   assign a0_mul_2x2_0 = a0x1; 
   assign a0_mul_2x2_1 = MASK1 ^ MASK2;
   assign a0_mul_2x3_0 = a0x2 ^ a0x7; 
   assign a0_mul_2x3_1 = MASK1;
   assign a0_mul_2x4_0 = a0x3 ^ a0x7; 
   assign a0_mul_2x4_1 = MASK1 ^ MASK2;
   assign a0_mul_2x5_0 = a0x4; 
   assign a0_mul_2x5_1 = MASK1;
   assign a0_mul_2x6_0 = a0x5; 
   assign a0_mul_2x6_1 = MASK2;
   assign a0_mul_2x7_0 = a0x6; 
   assign a0_mul_2x7_1 = MASK1;
   assign ha1x0_0 = a1x0^ MASK1; 
   assign ha1x0_1 = MASK1 ^ MASK2;
   assign a1_mul_2x0_0 = a1x7; 
   assign a1_mul_2x0_1 = MASK2;
   assign a1_mul_2x1_0 = ha1x0_0 ^ a1x7; 
   assign a1_mul_2x1_1 = MASK1;
   assign a1_mul_2x2_0 = a1x1; 
   assign a1_mul_2x2_1 = MASK1 ^ MASK2;
   assign a1_mul_2x3_0 = a1x2^ a1x7; 
   assign a1_mul_2x3_1 = MASK1;
   assign a1_mul_2x4_0 = a1x3^ a1x7; 
   assign a1_mul_2x4_1 = MASK1 ^ MASK2;
   assign a1_mul_2x5_0 = a1x4; 
   assign a1_mul_2x5_1 = MASK1;
   assign a1_mul_2x6_0 = a1x5; 
   assign a1_mul_2x6_1 = MASK2;
   assign a1_mul_2x7_0 = a1x6; 
   assign a1_mul_2x7_1 = MASK1;
   assign ha2x0_0 = a2x0 ^ MASK1; 
   assign ha2x0_1 = MASK1 ^ MASK2;
   assign a2_mul_2x0_0 = a2x7; 
   assign a2_mul_2x0_1 = MASK2;
   assign a2_mul_2x1_0 = ha2x0_0 ^ a2x7; 
   assign a2_mul_2x1_1 = MASK1;
   assign a2_mul_2x2_0 = a2x1; 
   assign a2_mul_2x2_1 = MASK1 ^ MASK2;
   assign a2_mul_2x3_0 = a2x2 ^ a2x7; 
   assign a2_mul_2x3_1 = MASK1;
   assign a2_mul_2x4_0 = a2x3 ^ a2x7; 
   assign a2_mul_2x4_1 = MASK1 ^ MASK2;
   assign a2_mul_2x5_0 = a2x4; 
   assign a2_mul_2x5_1 = MASK1;
   assign a2_mul_2x6_0 = a2x5; 
   assign a2_mul_2x6_1 = MASK2;
   assign a2_mul_2x7_0 = a2x6; 
   assign a2_mul_2x7_1 = MASK1;
   assign ha3x0_0 = a3x0 ^ MASK1; 
   assign ha3x0_1 = MASK1 ^ MASK2;
   assign a3_mul_2x0_0 = a3x7; 
   assign a3_mul_2x0_1 = MASK2;
   assign a3_mul_2x1_0 = ha3x0_0 ^ a3x7; 
   assign a3_mul_2x1_1 = MASK1;
   assign a3_mul_2x2_0 = a3x1; 
   assign a3_mul_2x2_1 = MASK1 ^ MASK2;
   assign a3_mul_2x3_0 = a3x2 ^ a3x7; 
   assign a3_mul_2x3_1 = MASK1;
   assign a3_mul_2x4_0 = a3x3 ^ a3x7; 
   assign a3_mul_2x4_1 = MASK1 ^ MASK2;
   assign a3_mul_2x5_0 = a3x4; 
   assign a3_mul_2x5_1 = MASK1;
   assign a3_mul_2x6_0 = a3x5; 
   assign a3_mul_2x6_1 = MASK2;
   assign a3_mul_2x7_0 = a3x6; 
   assign a3_mul_2x7_1 = MASK1;
   assign ha0_mul_2x0_0 = a0_mul_2x0_0 ^ MASK1; 
   assign ha0_mul_2x0_1 = MASK1 ^ MASK2;
   assign ha0_mul_2x2_0 = a0_mul_2x2_0 ^ MASK1; 
   assign ha0_mul_2x2_1 = MASK2;
   assign ha0_mul_2x3_0 = a0_mul_2x3_0 ^ MASK2; 
   assign ha0_mul_2x3_1 = MASK1 ^ MASK2;
   assign a0_mul_3x0_0 = ha0_mul_2x0_0 ^ a0x0; 
   assign a0_mul_3x0_1 = MASK1;
   assign a0_mul_3x1_0 = a0_mul_2x1_0 ^ a0x1; 
   assign a0_mul_3x1_1 = MASK2;
   assign a0_mul_3x2_0 = ha0_mul_2x2_0 ^ a0x2; 
   assign a0_mul_3x2_1 = MASK1;
   assign a0_mul_3x3_0 = ha0_mul_2x3_0 ^ a0x3; 
   assign a0_mul_3x3_1 = MASK2;
   assign a0_mul_3x4_0 = a0_mul_2x4_0 ^ a0x4; 
   assign a0_mul_3x4_1 = MASK2;
   assign a0_mul_3x5_0 = a0_mul_2x5_0 ^ a0x5; 
   assign a0_mul_3x5_1 = MASK1 ^ MASK2;
   assign a0_mul_3x6_0 = a0_mul_2x6_0 ^ a0x6; 
   assign a0_mul_3x6_1 = MASK1 ^ MASK2;
   assign a0_mul_3x7_0 = a0_mul_2x7_0 ^ a0x7; 
   assign a0_mul_3x7_1 = MASK1 ^ MASK2;
   assign ha1_mul_2x0_0 = a1_mul_2x0_0 ^ MASK1; 
   assign ha1_mul_2x0_1 = MASK1 ^ MASK2;
   assign ha1_mul_2x2_0 = a1_mul_2x2_0 ^ MASK1; 
   assign ha1_mul_2x2_1 = MASK2;
   assign ha1_mul_2x3_0 = a1_mul_2x3_0 ^ MASK2; 
   assign ha1_mul_2x3_1 = MASK1 ^ MASK2;
   assign a1_mul_3x0_0 = ha1_mul_2x0_0 ^ a1x0; 
   assign a1_mul_3x0_1 = MASK1;
   assign a1_mul_3x1_0 = a1_mul_2x1_0 ^ a1x1; 
   assign a1_mul_3x1_1 = MASK2;
   assign a1_mul_3x2_0 = ha1_mul_2x2_0 ^ a1x2; 
   assign a1_mul_3x2_1 = MASK1;
   assign a1_mul_3x3_0 = ha1_mul_2x3_0 ^ a1x3; 
   assign a1_mul_3x3_1 = MASK2;
   assign a1_mul_3x4_0 = a1_mul_2x4_0 ^ a1x4; 
   assign a1_mul_3x4_1 = MASK2;
   assign a1_mul_3x5_0 = a1_mul_2x5_0 ^ a1x5; 
   assign a1_mul_3x5_1 = MASK1 ^ MASK2;
   assign a1_mul_3x6_0 = a1_mul_2x6_0 ^ a1x6; 
   assign a1_mul_3x6_1 = MASK1 ^ MASK2;
   assign a1_mul_3x7_0 = a1_mul_2x7_0 ^ a1x7; 
   assign a1_mul_3x7_1 = MASK1 ^ MASK2;
   assign ha2_mul_2x0_0 = a2_mul_2x0_0 ^ MASK1; 
   assign ha2_mul_2x0_1 = MASK1 ^ MASK2;
   assign ha2_mul_2x2_0 = a2_mul_2x2_0 ^ MASK1; 
   assign ha2_mul_2x2_1 = MASK2;
   assign ha2_mul_2x3_0 = a2_mul_2x3_0 ^ MASK2; 
   assign ha2_mul_2x3_1 = MASK1 ^ MASK2;
   assign a2_mul_3x0_0 = ha2_mul_2x0_0 ^ a2x0; 
   assign a2_mul_3x0_1 = MASK1;
   assign a2_mul_3x1_0 = a2_mul_2x1_0 ^ a2x1; 
   assign a2_mul_3x1_1 = MASK2;
   assign a2_mul_3x2_0 = ha2_mul_2x2_0 ^ a2x2; 
   assign a2_mul_3x2_1 = MASK1;
   assign a2_mul_3x3_0 = ha2_mul_2x3_0 ^ a2x3; 
   assign a2_mul_3x3_1 = MASK2;
   assign a2_mul_3x4_0 = a2_mul_2x4_0 ^ a2x4; 
   assign a2_mul_3x4_1 = MASK2;
   assign a2_mul_3x5_0 = a2_mul_2x5_0 ^ a2x5; 
   assign a2_mul_3x5_1 = MASK1 ^ MASK2;
   assign a2_mul_3x6_0 = a2_mul_2x6_0 ^ a2x6; 
   assign a2_mul_3x6_1 = MASK1 ^ MASK2;
   assign a2_mul_3x7_0 = a2_mul_2x7_0 ^ a2x7; 
   assign a2_mul_3x7_1 = MASK1 ^ MASK2;
   assign ha3_mul_2x0_0 = a3_mul_2x0_0 ^ MASK1; 
   assign ha3_mul_2x0_1 = MASK1 ^ MASK2;
   assign ha3_mul_2x2_0 = a3_mul_2x2_0 ^ MASK1; 
   assign ha3_mul_2x2_1 = MASK2;
   assign ha3_mul_2x3_0 = a3_mul_2x3_0 ^ MASK2; 
   assign ha3_mul_2x3_1 = MASK1 ^ MASK2;
   assign a3_mul_3x0_0 = ha3_mul_2x0_0 ^ a3x0; 
   assign a3_mul_3x0_1 = MASK1;
   assign a3_mul_3x1_0 = a3_mul_2x1_0 ^ a3x1; 
   assign a3_mul_3x1_1 = MASK2;
   assign a3_mul_3x2_0 = ha3_mul_2x2_0 ^ a3x2; 
   assign a3_mul_3x2_1 = MASK1;
   assign a3_mul_3x3_0 = ha3_mul_2x3_0 ^ a3x3; 
   assign a3_mul_3x3_1 = MASK2;
   assign a3_mul_3x4_0 = a3_mul_2x4_0 ^ a3x4; 
   assign a3_mul_3x4_1 = MASK2;
   assign a3_mul_3x5_0 = a3_mul_2x5_0 ^ a3x5; 
   assign a3_mul_3x5_1 = MASK1 ^ MASK2;
   assign a3_mul_3x6_0 = a3_mul_2x6_0 ^ a3x6; 
   assign a3_mul_3x6_1 = MASK1 ^ MASK2;
   assign a3_mul_3x7_0 = a3_mul_2x7_0 ^ a3x7; 
   assign a3_mul_3x7_1 = MASK1 ^ MASK2;
   assign Ab0x0_0 = a0_mul_2x0_0 ^ a1_mul_3x0_0; 
   assign Ab0x0_1 = MASK1 ^ MASK2;
   assign Ab0x1_0 = a0_mul_2x1_0 ^ a1_mul_3x1_0; 
   assign Ab0x1_1 = MASK1 ^ MASK2;
   assign Ab0x2_0 = a0_mul_2x2_0 ^ a1_mul_3x2_0; 
   assign Ab0x2_1 = MASK2;
   assign Ab0x3_0 = a0_mul_2x3_0 ^ a1_mul_3x3_0; 
   assign Ab0x3_1 = MASK1 ^ MASK2;
   assign Ab0x4_0 = a0_mul_2x4_0 ^ a1_mul_3x4_0; 
   assign Ab0x4_1 = MASK1;
   assign Ab0x5_0 = a0_mul_2x5_0 ^ a1_mul_3x5_0; 
   assign Ab0x5_1 = MASK2;
   assign Ab0x6_0 = a0_mul_2x6_0 ^ a1_mul_3x6_0; 
   assign Ab0x6_1 = MASK1;
   assign Ab0x7_0 = a0_mul_2x7_0 ^ a1_mul_3x7_0; 
   assign Ab0x7_1 = MASK2;
   assign ha3x1_0 = a3x1 ^ MASK1; 
   assign ha3x1_1 = MASK2;
   assign ha3x2_0 = a3x2 ^ MASK1; 
   assign ha3x2_1 = MASK2;
   assign ha3x3_0 = a3x3 ^ MASK2; 
   assign ha3x3_1 = MASK1 ^ MASK2;
   assign ha3x4_0 = a3x4 ^ MASK2; 
   assign ha3x4_1 = MASK1 ^ MASK2;
   assign ha3x5_0 = a3x5 ^ MASK1; 
   assign ha3x5_1 = MASK1 ^ MASK2;
   assign ha3x6_0 = a3x6 ^ MASK2; 
   assign ha3x6_1 = MASK1 ^ MASK2;
   assign ha3x7_0 = a3x7 ^ MASK1; 
   assign ha3x7_1 = MASK1 ^ MASK2;
   assign Bb0x0_0 = ha2x0_0 ^ a3x0; 
   assign Bb0x0_1 = MASK1;
   assign Bb0x1_0 = a2x1 ^ ha3x1_0; 
   assign Bb0x1_1 = MASK1;
   assign Bb0x2_0 = a2x2 ^ ha3x2_0; 
   assign Bb0x2_1 = MASK1;
   assign Bb0x3_0 = a2x3 ^ ha3x3_0; 
   assign Bb0x3_1 = MASK2;
   assign Bb0x4_0 = a2x4 ^ ha3x4_0; 
   assign Bb0x4_1 = MASK2;
   assign Bb0x5_0 = a2x5 ^ ha3x5_0; 
   assign Bb0x5_1 = MASK1;
   assign Bb0x6_0 = a2x6 ^ ha3x6_0; 
   assign Bb0x6_1 = MASK2;
   assign Bb0x7_0 = a2x7^ ha3x7_0; 
   assign Bb0x7_1 = MASK1;
   assign b0x0 = Ab0x0_0 ^ Bb0x0_0; 
   assign hb0x1_0 = Ab0x1_0 ^ Bb0x1_0; 
   assign hb0x1_1 = MASK2;
   assign b0x1 = hb0x1_0 ^ MASK1; 
   assign hb0x2_0 = Ab0x2_0 ^ Bb0x2_0; 
   assign hb0x2_1 = MASK1 ^ MASK2;
   assign b0x2 = hb0x2_0; 
   assign b0x3 = Ab0x3_0 ^ Bb0x3_0; 
   assign hb0x4_0 = Ab0x4_0 ^ Bb0x4_0; 
   assign hb0x4_1 = MASK1 ^ MASK2;
   assign b0x4 = hb0x4_0 ^ MASK2; 
   assign hb0x5_0 = Ab0x5_0 ^ Bb0x5_0; 
   assign hb0x5_1 = MASK1 ^ MASK2;
   assign b0x5 = hb0x5_0 ^ MASK1; 
   assign hb0x6_0 = Ab0x6_0 ^ Bb0x6_0; 
   assign hb0x6_1 = MASK1 ^ MASK2;
   assign b0x6 = hb0x6_0 ^ MASK2; 
   assign hb0x7_0 = Ab0x7_0 ^ Bb0x7_0; 
   assign hb0x7_1 = MASK1 ^ MASK2;
   assign b0x7 = hb0x7_0 ^ MASK1; 
   assign Ab1x0_0 = ha0x0_0 ^ a1_mul_2x0_0; 
   assign Ab1x0_1 = MASK1;
   assign Ab1x1_0 = a0x1 ^ a1_mul_2x1_0; 
   assign Ab1x1_1 = MASK2;
   assign Ab1x2_0 = a0x2 ^ ha1_mul_2x2_0; 
   assign Ab1x2_1 = MASK1;
   assign Ab1x3_0 = a0x3^ ha1_mul_2x3_0; 
   assign Ab1x3_1 = MASK2;
   assign Ab1x4_0 = a0x4^ a1_mul_2x4_0; 
   assign Ab1x4_1 = MASK2;
   assign Ab1x5_0 = a0x5^ a1_mul_2x5_0; 
   assign Ab1x5_1 = MASK1 ^ MASK2;
   assign Ab1x6_0 = a0x6^ a1_mul_2x6_0; 
   assign Ab1x6_1 = MASK1 ^ MASK2;
   assign Ab1x7_0 = a0x7^ a1_mul_2x7_0; 
   assign Ab1x7_1 = MASK1 ^ MASK2;
   assign Bb1x0_0 = a2_mul_3x0_0 ^ a3x0; 
   assign Bb1x0_1 = MASK1 ^ MASK2;
   assign Bb1x1_0 = a2_mul_3x1_0 ^ a3x1; 
   assign Bb1x1_1 = MASK1;
   assign Bb1x2_0 = a2_mul_3x2_0 ^ a3x2; 
   assign Bb1x2_1 = MASK2;
   assign Bb1x3_0 = a2_mul_3x3_0 ^ a3x3; 
   assign Bb1x3_1 = MASK1 ^ MASK2;
   assign Bb1x4_0 = a2_mul_3x4_0 ^ a3x4; 
   assign Bb1x4_1 = MASK1 ^ MASK2;
   assign Bb1x5_0 = a2_mul_3x5_0 ^ a3x5; 
   assign Bb1x5_1 = MASK1;
   assign Bb1x6_0 = a2_mul_3x6_0 ^ a3x6; 
   assign Bb1x6_1 = MASK2;
   assign Bb1x7_0 = a2_mul_3x7_0 ^ a3x7; 
   assign Bb1x7_1 = MASK1;
   assign b1x0 = Ab1x0_0 ^ Bb1x0_0; 
   assign b1x1 = Ab1x1_0 ^ Bb1x1_0; 
   assign b1x2 = Ab1x2_0 ^ Bb1x2_0; 
   assign b1x3 = Ab1x3_0 ^ Bb1x3_0; 
   assign b1x4 = Ab1x4_0 ^ Bb1x4_0; 
   assign b1x5 = Ab1x5_0 ^ Bb1x5_0; 
   assign b1x6 = Ab1x6_0 ^ Bb1x6_0; 
   assign b1x7 = Ab1x7_0 ^ Bb1x7_0; 
   assign ha0x1_0 = a0x1 ^ MASK1; 
   assign ha0x1_1 = MASK2;
   assign ha0x2_0 = a0x2 ^ MASK1; 
   assign ha0x2_1 = MASK2;
   assign ha0x3_0 = a0x3^ MASK2; 
   assign ha0x3_1 = MASK1 ^ MASK2;
   assign ha0x4_0 = a0x4^ MASK2; 
   assign ha0x4_1 = MASK1 ^ MASK2;
   assign ha0x5_0 = a0x5^ MASK1; 
   assign ha0x5_1 = MASK1 ^ MASK2;
   assign ha0x6_0 = a0x6^ MASK2; 
   assign ha0x6_1 = MASK1 ^ MASK2;
   assign ha0x7_0 = a0x7^ MASK1; 
   assign ha0x7_1 = MASK1 ^ MASK2;
   assign Ab2x0_0 = ha0x0_0 ^ a1x0; 
   assign Ab2x0_1 = MASK1;
   assign Ab2x1_0 = ha0x1_0 ^ a1x1; 
   assign Ab2x1_1 = MASK1;
   assign Ab2x2_0 = ha0x2_0 ^ a1x2; 
   assign Ab2x2_1 = MASK1;
   assign Ab2x3_0 = ha0x3_0 ^ a1x3; 
   assign Ab2x3_1 = MASK2;
   assign Ab2x4_0 = ha0x4_0 ^ a1x4; 
   assign Ab2x4_1 = MASK2;
   assign Ab2x5_0 = ha0x5_0 ^ a1x5; 
   assign Ab2x5_1 = MASK1;
   assign Ab2x6_0 = ha0x6_0 ^ a1x6; 
   assign Ab2x6_1 = MASK2;
   assign Ab2x7_0 = ha0x7_0 ^ a1x7; 
   assign Ab2x7_1 = MASK1;
   assign Bb2x0_0 = a2_mul_2x0_0 ^ a3_mul_3x0_0; 
   assign Bb2x0_1 = MASK1 ^ MASK2;
   assign Bb2x1_0 = a2_mul_2x1_0 ^ a3_mul_3x1_0; 
   assign Bb2x1_1 = MASK1 ^ MASK2;
   assign Bb2x2_0 = a2_mul_2x2_0 ^ a3_mul_3x2_0; 
   assign Bb2x2_1 = MASK2;
   assign Bb2x3_0 = a2_mul_2x3_0 ^ a3_mul_3x3_0; 
   assign Bb2x3_1 = MASK1 ^ MASK2;
   assign Bb2x4_0 = a2_mul_2x4_0 ^ a3_mul_3x4_0; 
   assign Bb2x4_1 = MASK1;
   assign Bb2x5_0 = a2_mul_2x5_0 ^ a3_mul_3x5_0; 
   assign Bb2x5_1 = MASK2;
   assign Bb2x6_0 = a2_mul_2x6_0 ^ a3_mul_3x6_0; 
   assign Bb2x6_1 = MASK1;
   assign Bb2x7_0 = a2_mul_2x7_0 ^ a3_mul_3x7_0; 
   assign Bb2x7_1 = MASK2;
   assign b2x0 = Ab2x0_0 ^ Bb2x0_0; 
   assign hb2x1_0 = Ab2x1_0 ^ Bb2x1_0; 
   assign hb2x1_1 = MASK2;
   assign b2x1 = hb2x1_0 ^ MASK1; 
   assign b2x2 = Ab2x2_0 ^ Bb2x2_0; 
   assign b2x3 = Ab2x3_0 ^ Bb2x3_0; 
   assign hb2x4_0 = Ab2x4_0 ^ Bb2x4_0; 
   assign hb2x4_1 = MASK1 ^ MASK2;
   assign b2x4 = hb2x4_0 ^ MASK2; 
   assign hb2x5_0 = Ab2x5_0 ^ Bb2x5_0; 
   assign hb2x5_1 = MASK1 ^ MASK2;
   assign b2x5 = hb2x5_0 ^ MASK1; 
   assign hb2x6_0 = Ab2x6_0 ^ Bb2x6_0; 
   assign hb2x6_1 = MASK1 ^ MASK2;
   assign b2x6 = hb2x6_0 ^ MASK2; 
   assign hb2x7_0 = Ab2x7_0 ^ Bb2x7_0; 
   assign hb2x7_1 = MASK1 ^ MASK2;
   assign b2x7 = hb2x7_0 ^ MASK1; 
   assign Ab3x0_0 = a0_mul_3x0_0 ^ a1x0; 
   assign Ab3x0_1 = MASK1 ^ MASK2;
   assign Ab3x1_0 = a0_mul_3x1_0 ^ a1x1; 
   assign Ab3x1_1 = MASK1;             
   assign Ab3x2_0 = a0_mul_3x2_0 ^ a1x2; 
   assign Ab3x2_1 = MASK2;
   assign Ab3x3_0 = a0_mul_3x3_0 ^ a1x3; 
   assign Ab3x3_1 = MASK1 ^ MASK2;
   assign Ab3x4_0 = a0_mul_3x4_0 ^ a1x4; 
   assign Ab3x4_1 = MASK1 ^ MASK2;     
   assign Ab3x5_0 = a0_mul_3x5_0 ^ a1x5; 
   assign Ab3x5_1 = MASK1;
   assign Ab3x6_0 = a0_mul_3x6_0 ^ a1x6; 
   assign Ab3x6_1 = MASK2;
   assign Ab3x7_0 = a0_mul_3x7_0 ^ a1x7; 
   assign Ab3x7_1 = MASK1;
   assign Bb3x0_0 = ha2x0_0 ^ a3_mul_2x0_0; 
   assign Bb3x0_1 = MASK1;
   assign Bb3x1_0 = a2x1 ^ a3_mul_2x1_0; 
   assign Bb3x1_1 = MASK2;
   assign Bb3x2_0 = a2x2 ^ ha3_mul_2x2_0; 
   assign Bb3x2_1 = MASK1;
   assign Bb3x3_0 = a2x3 ^ ha3_mul_2x3_0; 
   assign Bb3x3_1 = MASK2;
   assign Bb3x4_0 = a2x4 ^ a3_mul_2x4_0; 
   assign Bb3x4_1 = MASK2;
   assign Bb3x5_0 = a2x5 ^ a3_mul_2x5_0; 
   assign Bb3x5_1 = MASK1 ^ MASK2;
   assign Bb3x6_0 = a2x6 ^ a3_mul_2x6_0; 
   assign Bb3x6_1 = MASK1 ^ MASK2;
   assign Bb3x7_0 = a2x7^ a3_mul_2x7_0; 
   assign Bb3x7_1 = MASK1 ^ MASK2;
   assign b3x0 = Ab3x0_0 ^ Bb3x0_0; 
   assign b3x1 = Ab3x1_0 ^ Bb3x1_0; 
   assign b3x2 = Ab3x2_0 ^ Bb3x2_0; 
   assign b3x3 = Ab3x3_0 ^ Bb3x3_0; 
   assign b3x4 = Ab3x4_0 ^ Bb3x4_0; 
   assign b3x5 = Ab3x5_0 ^ Bb3x5_0; 
   assign b3x6 = Ab3x6_0 ^ Bb3x6_0; 
   assign b3x7 = Ab3x7_0 ^ Bb3x7_0; 

endmodule // mixcolumns